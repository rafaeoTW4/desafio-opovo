<svg width="29" height="18" viewBox="0 0 29 18" fill="none" xmlns="http://www.w3.org/2000/svg">
<path d="M2 2.75L14.5 15.25L27 2.75" stroke="#1F6482" stroke-width="4" stroke-linecap="round" stroke-linejoin="round"/>
</svg>
